//2252429������
`timescale 1ns / 1ps
//cpu31��������ģ��
module cpu31_tb();
//---------------------------------------------------------------   
    //�����ڲ�����
    reg clk;                    //ʱ���ź�
    reg rst;                    //��λ�ź�
    wire [31:0] inst;           //ִ�е�ָ��
    wire [31:0] pc;             //��һ��ָ��ĵ�ַ
//---------------------------------------------------------------   
//cpuʵ����
sccomp_dataflow cpu31_inst(
    .clk_in(clk),
    .reset(rst),
    .inst(inst),
    .pc(pc)
);
//---------------------------------------------------------------   
initial 
    begin
    clk = 0;
    rst = 1;
    //wait for gloabal rest to finish
    #50
    rst = 0;
    end
//---------------------------------------------------------------   
//����ʱ��
    always #50 clk =~clk;
//---------------------------------------------------------------   
endmodule
